/////////////////////////////////////////////////////////////////////////////////////
// Copyright 2019 seabeam@yahoo.com - Licensed under the Apache License, Version 2.0
// For more information, see LICENCE in the main folder
/////////////////////////////////////////////////////////////////////////////////////
`ifndef YUU_CLOCK_DEFINES_SVH
`define YUU_CLOCK_DEFINES_SVH

  `ifndef YUU_CLOCK_MAX_DIVIDE
  `define YUU_CLOCK_MAX_DIVIDE  16
  `endif

  `ifndef YUU_CLOCK_MAX_MULTI
  `define YUU_CLOCK_MAX_MULTI   16
  `endif
  
`endif
